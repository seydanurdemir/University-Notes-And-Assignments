magic
tech scmos
timestamp 1606509372
<< ntransistor >>
rect 6 0 8 4
rect 16 0 18 4
<< ptransistor >>
rect 6 16 8 20
rect 16 16 18 20
<< ndiffusion >>
rect 4 0 6 4
rect 8 0 10 4
rect 14 0 16 4
rect 18 0 20 4
<< pdiffusion >>
rect 4 16 6 20
rect 8 16 16 20
rect 18 16 20 20
<< ndcontact >>
rect 0 0 4 4
rect 10 0 14 4
rect 20 0 24 4
<< pdcontact >>
rect 0 16 4 20
rect 20 16 24 20
<< polysilicon >>
rect 6 20 8 23
rect 16 20 18 23
rect 6 4 8 16
rect 16 4 18 16
rect 6 -3 8 0
rect 16 -3 18 0
<< metal1 >>
rect 0 20 4 24
rect 20 12 24 16
rect 10 8 24 12
rect 10 4 14 8
rect 0 -4 4 0
rect 20 -4 24 0
rect 0 -8 24 -4
<< labels >>
rlabel pdcontact 2 18 2 18 1 VDD
rlabel ndcontact 2 2 2 2 1 GND
rlabel polysilicon 7 14 7 14 1 A
rlabel polysilicon 17 14 17 14 1 B
rlabel metal1 22 14 22 14 1 Z
<< end >>
