magic
tech scmos
timestamp 1606508494
<< ntransistor >>
rect 6 0 8 4
rect 16 0 18 4
<< ptransistor >>
rect 6 16 8 20
rect 16 16 18 20
<< ndiffusion >>
rect 4 0 6 4
rect 8 0 16 4
rect 18 0 20 4
<< pdiffusion >>
rect 4 16 6 20
rect 8 16 10 20
rect 14 16 16 20
rect 18 16 20 20
<< ndcontact >>
rect 0 0 4 4
rect 20 0 24 4
<< pdcontact >>
rect 0 16 4 20
rect 10 16 14 20
rect 20 16 24 20
<< polysilicon >>
rect 6 20 8 23
rect 16 20 18 23
rect 6 4 8 16
rect 16 4 18 16
rect 6 -3 8 0
rect 16 -3 18 0
<< metal1 >>
rect 0 24 24 27
rect 0 20 4 24
rect 20 20 24 24
rect 10 12 14 16
rect 10 8 24 12
rect 20 4 24 8
rect 0 -4 4 0
<< labels >>
rlabel ndcontact 2 2 2 2 1 GND
rlabel pdcontact 2 18 2 18 1 VDD
rlabel metal1 22 6 22 6 1 Z
rlabel polysilicon 17 6 17 6 1 B
rlabel polysilicon 7 6 7 6 1 A
<< end >>
